//name : main_0
//input : input_eth_in:16
//output : output_eth_out:16
//output : output_rs232_out:16
//source_file : /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_eth_in,input_eth_in_stb,output_eth_out_ack,output_rs232_out_ack,clk,rst,output_eth_out,output_rs232_out,output_eth_out_stb,output_rs232_out_stb,input_eth_in_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_eth_in;
  input input_eth_in_stb;
  input output_eth_out_ack;
  input output_rs232_out_ack;
  input clk;
  input rst;
  output [31:0] output_eth_out;
  output [31:0] output_rs232_out;
  output output_eth_out_stb;
  output output_rs232_out_stb;
  output input_eth_in_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_eth_out_stb;
  reg [31:0] s_output_rs232_out_stb;
  reg [31:0] s_output_eth_out;
  reg [31:0] s_output_rs232_out;
  reg [31:0] s_input_eth_in_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [925:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': False, 'op': 'add'}
  // 7 {'literal': False, 'op': 'greater'}
  // 8 {'literal': True, 'op': 'jmp_if_false'}
  // 9 {'literal': False, 'op': 'shift_left'}
  // 10 {'literal': False, 'op': 'subtract'}
  // 11 {'literal': True, 'op': 'goto'}
  // 12 {'literal': False, 'op': 'return'}
  // 13 {'literal': False, 'op': 'write'}
  // 14 {'literal': False, 'op': 'read'}
  // 15 {'literal': False, 'op': 'unsigned_shift_right'}
  // 16 {'literal': False, 'op': 'equal'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd43};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'a': 3, 'literal': 43, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7 {'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7 {'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 7, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6 {'literal': 2, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 6, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd3};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd5};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1 {'literal': 5, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 1, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd67};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 67, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 8, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd104};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 104, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd9};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 9, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd105};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 105, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 10, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd112};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 112, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd11};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 11, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd115};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 115, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd12};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 12, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd32};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 32, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd13};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 13, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd105};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 105, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd14};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 14, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd109};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 109, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd15};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 15, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd97};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 97, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd16};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 16, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd103};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 103, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd17};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 17, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd18};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 18, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd32};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 32, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd19};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 19, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd112};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 112, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd20};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 20, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd114};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 114, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd21};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 21, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd111};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 111, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd22};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 22, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd99};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 99, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd23};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 23, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd24};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 24, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd115};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 115, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd25};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 25, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd115};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 115, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd26};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 26, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd105};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 105, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd27};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 27, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd110};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 110, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd28};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 28, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd103};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 103, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd29};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 29, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd32};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 32, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd30};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 30, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd31};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 31, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd120};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 120, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd32};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 32, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd97};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 97, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd33};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 33, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd109};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 109, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd34};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 34, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd112};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 112, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd35};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 35, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd108};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 108, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd36};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 36, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd37};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 37, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 10, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd38};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 38, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd39};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 39, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3 {'literal': 1029, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd40};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3 {'literal': 40, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 3, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5 {'literal': 41, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 5, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd515};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2 {'literal': 515, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd42};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2 {'literal': 42, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 2, 'op': 'store'}
    instructions[120] = {5'd1, 4'd7, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'addl'}
    instructions[121] = {5'd1, 4'd4, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'addl'}
    instructions[122] = {5'd3, 4'd6, 4'd0, 16'd124};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'z': 6, 'label': 124, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'call'}
    instructions[123] = {5'd4, 4'd0, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72 {'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 72, 'op': 'stop'}
    instructions[124] = {5'd1, 4'd3, 4'd3, 16'd132135};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25 {'a': 3, 'literal': 132135, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25, 'op': 'addl'}
    instructions[125] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39 {'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39, 'op': 'literal'}
    instructions[126] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39, 'op': 'addl'}
    instructions[127] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39, 'op': 'load'}
    instructions[128] = {5'd0, 4'd2, 4'd0, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39 {'literal': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39, 'op': 'literal'}
    instructions[129] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 39, 'op': 'store'}
    instructions[130] = {5'd2, 4'd0, 4'd3, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[131] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[132] = {5'd2, 4'd0, 4'd3, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[133] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[134] = {5'd0, 4'd8, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'literal': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'literal'}
    instructions[135] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'store'}
    instructions[136] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[137] = {5'd1, 4'd7, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[138] = {5'd1, 4'd4, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[139] = {5'd3, 4'd6, 4'd0, 16'd438};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'z': 6, 'label': 438, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'call'}
    instructions[140] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[141] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[142] = {5'd5, 4'd7, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'load'}
    instructions[143] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[144] = {5'd5, 4'd6, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'z': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'load'}
    instructions[145] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 41, 'op': 'addl'}
    instructions[146] = {5'd1, 4'd8, 4'd4, 16'd131075};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 4, 'literal': 131075, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'addl'}
    instructions[147] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'store'}
    instructions[148] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'addl'}
    instructions[149] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'literal'}
    instructions[150] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[151] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'load'}
    instructions[152] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'add'}
    instructions[153] = {5'd1, 4'd2, 4'd4, 16'd132099};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 4, 'literal': 132099, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'addl'}
    instructions[154] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 43, 'op': 'store'}
    instructions[155] = {5'd1, 4'd8, 4'd4, 16'd131331};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 4, 'literal': 131331, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'addl'}
    instructions[156] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'store'}
    instructions[157] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'addl'}
    instructions[158] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'literal'}
    instructions[159] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[160] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'load'}
    instructions[161] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'add'}
    instructions[162] = {5'd1, 4'd2, 4'd4, 16'd132100};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 4, 'literal': 132100, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'addl'}
    instructions[163] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 44, 'op': 'store'}
    instructions[164] = {5'd1, 4'd8, 4'd4, 16'd131587};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 4, 'literal': 131587, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'addl'}
    instructions[165] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'store'}
    instructions[166] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'addl'}
    instructions[167] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'literal'}
    instructions[168] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[169] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'load'}
    instructions[170] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'add'}
    instructions[171] = {5'd1, 4'd2, 4'd4, 16'd132101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 4, 'literal': 132101, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'addl'}
    instructions[172] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 45, 'op': 'store'}
    instructions[173] = {5'd1, 4'd8, 4'd4, 16'd132100};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50 {'a': 4, 'literal': 132100, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50, 'op': 'addl'}
    instructions[174] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50, 'op': 'addl'}
    instructions[175] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50, 'op': 'load'}
    instructions[176] = {5'd1, 4'd2, 4'd4, 16'd132101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50 {'a': 4, 'literal': 132101, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50, 'op': 'addl'}
    instructions[177] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 50, 'op': 'store'}
    instructions[178] = {5'd1, 4'd8, 4'd4, 16'd132099};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51 {'a': 4, 'literal': 132099, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51, 'op': 'addl'}
    instructions[179] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51, 'op': 'addl'}
    instructions[180] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51, 'op': 'load'}
    instructions[181] = {5'd1, 4'd2, 4'd4, 16'd132100};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51 {'a': 4, 'literal': 132100, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51, 'op': 'addl'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 51, 'op': 'store'}
    instructions[183] = {5'd2, 4'd0, 4'd3, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'store'}
    instructions[184] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[185] = {5'd2, 4'd0, 4'd3, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'store'}
    instructions[186] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[187] = {5'd1, 4'd8, 4'd4, 16'd132099};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 4, 'literal': 132099, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[188] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[189] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'load'}
    instructions[190] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'store'}
    instructions[191] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[192] = {5'd1, 4'd7, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[193] = {5'd1, 4'd4, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[194] = {5'd3, 4'd6, 4'd0, 16'd529};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'z': 6, 'label': 529, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'call'}
    instructions[195] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[196] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[197] = {5'd5, 4'd7, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'load'}
    instructions[198] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[199] = {5'd5, 4'd6, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 3, 'z': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'load'}
    instructions[200] = {5'd0, 4'd2, 4'd0, 16'd4};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'literal': 4, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'literal'}
    instructions[201] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'load'}
    instructions[202] = {5'd1, 4'd2, 4'd4, 16'd132102};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 4, 'literal': 132102, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'addl'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 52, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'literal'}
    instructions[205] = {5'd1, 4'd2, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 4, 'literal': 131072, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'store'}
    instructions[207] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[208] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[209] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[210] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'store'}
    instructions[211] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[212] = {5'd0, 4'd8, 4'd0, 16'd256};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'literal': 256, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'literal'}
    instructions[213] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[214] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[215] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'greater'}
    instructions[216] = {5'd8, 4'd0, 4'd8, 16'd413};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'label': 413, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'jmp_if_false'}
    instructions[217] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'store'}
    instructions[219] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[220] = {5'd1, 4'd8, 4'd4, 16'd132100};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 4, 'literal': 132100, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[221] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[222] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'load'}
    instructions[223] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'store'}
    instructions[224] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[225] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[226] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[227] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'load'}
    instructions[228] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[229] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'load'}
    instructions[230] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'add'}
    instructions[231] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[232] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'load'}
    instructions[233] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[234] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'load'}
    instructions[235] = {5'd9, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'shift_left'}
    instructions[236] = {5'd1, 4'd2, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 4, 'literal': 131074, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'addl'}
    instructions[237] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 55, 'op': 'store'}
    instructions[238] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'literal'}
    instructions[239] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'store'}
    instructions[240] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'addl'}
    instructions[241] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'addl'}
    instructions[242] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'addl'}
    instructions[243] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'load'}
    instructions[244] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[245] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'load'}
    instructions[246] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'greater'}
    instructions[247] = {5'd8, 4'd0, 4'd8, 16'd307};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'a': 8, 'label': 307, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'jmp_if_false'}
    instructions[248] = {5'd1, 4'd8, 4'd4, 16'd132099};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 4, 'literal': 132099, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[249] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[250] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[251] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'store'}
    instructions[252] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[253] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'literal'}
    instructions[254] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'store'}
    instructions[255] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[256] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[257] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[258] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[259] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[260] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[261] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'subtract'}
    instructions[262] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[263] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[264] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'add'}
    instructions[265] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[266] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[267] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'store'}
    instructions[268] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[269] = {5'd1, 4'd8, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 4, 'literal': 131074, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[270] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[271] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[272] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[273] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'load'}
    instructions[274] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'subtract'}
    instructions[275] = {5'd1, 4'd2, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 4, 'literal': 131074, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'addl'}
    instructions[276] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 57, 'op': 'store'}
    instructions[277] = {5'd1, 4'd8, 4'd4, 16'd132101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 4, 'literal': 132101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[278] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[279] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[280] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'store'}
    instructions[281] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'literal'}
    instructions[283] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'store'}
    instructions[284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[285] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[286] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[287] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[288] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[289] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[290] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'subtract'}
    instructions[291] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[292] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[293] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'add'}
    instructions[294] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[295] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[296] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'store'}
    instructions[297] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[298] = {5'd1, 4'd8, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 4, 'literal': 131074, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[299] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[300] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[301] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[302] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'load'}
    instructions[303] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'subtract'}
    instructions[304] = {5'd1, 4'd2, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 4, 'literal': 131074, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'addl'}
    instructions[305] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 58, 'op': 'store'}
    instructions[306] = {5'd11, 4'd0, 4'd0, 16'd307};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56 {'label': 307, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 56, 'op': 'goto'}
    instructions[307] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'addl'}
    instructions[308] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'addl'}
    instructions[309] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'load'}
    instructions[310] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'store'}
    instructions[311] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'addl'}
    instructions[312] = {5'd0, 4'd8, 4'd0, 16'd255};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'literal': 255, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'literal'}
    instructions[313] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[314] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'load'}
    instructions[315] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'greater'}
    instructions[316] = {5'd8, 4'd0, 4'd8, 16'd376};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'a': 8, 'label': 376, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'jmp_if_false'}
    instructions[317] = {5'd1, 4'd8, 4'd4, 16'd132101};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 4, 'literal': 132101, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[318] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[319] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[320] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'store'}
    instructions[321] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[322] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'literal'}
    instructions[323] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'store'}
    instructions[324] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[325] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[326] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[327] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[328] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[329] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[330] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'add'}
    instructions[331] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[332] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[333] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'add'}
    instructions[334] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[335] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[336] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'store'}
    instructions[337] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[338] = {5'd1, 4'd8, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 4, 'literal': 131074, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[339] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[340] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[341] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[342] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'load'}
    instructions[343] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'subtract'}
    instructions[344] = {5'd1, 4'd2, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 4, 'literal': 131074, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'addl'}
    instructions[345] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 61, 'op': 'store'}
    instructions[346] = {5'd1, 4'd8, 4'd4, 16'd132099};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 4, 'literal': 132099, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[347] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[348] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[349] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'store'}
    instructions[350] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[351] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'literal'}
    instructions[352] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'store'}
    instructions[353] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[354] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[355] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[356] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[357] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[358] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[359] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'add'}
    instructions[360] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[361] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[362] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'add'}
    instructions[363] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[364] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[365] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'store'}
    instructions[366] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[367] = {5'd1, 4'd8, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 4, 'literal': 131074, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[368] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[369] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[370] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[371] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'load'}
    instructions[372] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'subtract'}
    instructions[373] = {5'd1, 4'd2, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 4, 'literal': 131074, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'addl'}
    instructions[374] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 62, 'op': 'store'}
    instructions[375] = {5'd11, 4'd0, 4'd0, 16'd376};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60 {'label': 376, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 60, 'op': 'goto'}
    instructions[376] = {5'd1, 4'd8, 4'd4, 16'd131074};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 4, 'literal': 131074, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[377] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[378] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'load'}
    instructions[379] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'store'}
    instructions[380] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[381] = {5'd1, 4'd8, 4'd4, 16'd131843};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 4, 'literal': 131843, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[382] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'store'}
    instructions[383] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[384] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[385] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[386] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'load'}
    instructions[387] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[388] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'load'}
    instructions[389] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'add'}
    instructions[390] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'addl'}
    instructions[391] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[392] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'load'}
    instructions[393] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 64, 'op': 'store'}
    instructions[394] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[395] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[396] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[397] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'store'}
    instructions[398] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[399] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'literal'}
    instructions[400] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'store'}
    instructions[401] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[402] = {5'd1, 4'd8, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 4, 'literal': 131072, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[403] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[404] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[405] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[406] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[407] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'add'}
    instructions[408] = {5'd1, 4'd2, 4'd4, 16'd131072};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 4, 'literal': 131072, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'addl'}
    instructions[409] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'store'}
    instructions[410] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[411] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'load'}
    instructions[412] = {5'd11, 4'd0, 4'd0, 16'd207};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54 {'label': 207, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 54, 'op': 'goto'}
    instructions[413] = {5'd2, 4'd0, 4'd3, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'store'}
    instructions[414] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[415] = {5'd2, 4'd0, 4'd3, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'store'}
    instructions[416] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[417] = {5'd1, 4'd8, 4'd4, 16'd131843};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 4, 'literal': 131843, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[418] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'store'}
    instructions[419] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[420] = {5'd1, 4'd8, 4'd4, 16'd132102};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 4, 'literal': 132102, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[421] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[422] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'load'}
    instructions[423] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'store'}
    instructions[424] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[425] = {5'd1, 4'd7, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[426] = {5'd1, 4'd4, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[427] = {5'd3, 4'd6, 4'd0, 16'd739};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'z': 6, 'label': 739, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'call'}
    instructions[428] = {5'd1, 4'd3, 4'd3, -16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[429] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[430] = {5'd5, 4'd7, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'z': 7, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'load'}
    instructions[431] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[432] = {5'd5, 4'd6, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'z': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'load'}
    instructions[433] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 67, 'op': 'addl'}
    instructions[434] = {5'd11, 4'd0, 4'd0, 16'd173};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 46 {'label': 173, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 46, 'op': 'goto'}
    instructions[435] = {5'd1, 4'd3, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25, 'op': 'addl'}
    instructions[436] = {5'd1, 4'd4, 4'd7, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25, 'op': 'addl'}
    instructions[437] = {5'd12, 4'd0, 4'd6, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25 {'a': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/application.c : 25, 'op': 'return'}
    instructions[438] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[439] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[440] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[441] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[442] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[443] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[444] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[445] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[446] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[447] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[448] = {5'd0, 4'd8, 4'd0, 16'd3};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[449] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[450] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[451] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[452] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[453] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[454] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[455] = {5'd3, 4'd6, 4'd0, 16'd465};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 465, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[456] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[457] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[458] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[459] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[460] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[461] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[462] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[463] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[464] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[465] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[466] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[467] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[468] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[469] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[470] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[471] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[472] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[473] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[474] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[475] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[476] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[477] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[478] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[479] = {5'd6, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[480] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[481] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[482] = {5'd8, 4'd0, 4'd8, 16'd524};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 524, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[483] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[484] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[485] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[486] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[487] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[488] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[489] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[490] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[491] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[492] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[493] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[494] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[495] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[496] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[497] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[498] = {5'd6, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[499] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[500] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[501] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[502] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[503] = {5'd13, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[504] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[505] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[506] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[507] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[508] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[509] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[510] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[511] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[512] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[513] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[514] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[515] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[516] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[517] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[518] = {5'd6, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[519] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[520] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[521] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[522] = {5'd5, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[523] = {5'd11, 4'd0, 4'd0, 16'd525};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 525, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[524] = {5'd11, 4'd0, 4'd0, 16'd526};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 526, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[525] = {5'd11, 4'd0, 4'd0, 16'd469};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 469, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[526] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[527] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[528] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[529] = {5'd1, 4'd3, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 7 {'a': 3, 'literal': 8, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 7, 'op': 'addl'}
    instructions[530] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'literal'}
    instructions[531] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'addl'}
    instructions[532] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'load'}
    instructions[533] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'read'}
    instructions[534] = {5'd1, 4'd2, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'addl'}
    instructions[535] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 13, 'op': 'store'}
    instructions[536] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'literal'}
    instructions[537] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'addl'}
    instructions[538] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'load'}
    instructions[539] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'read'}
    instructions[540] = {5'd1, 4'd2, 4'd4, 16'd4};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'addl'}
    instructions[541] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 14, 'op': 'store'}
    instructions[542] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'literal'}
    instructions[543] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'addl'}
    instructions[544] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'load'}
    instructions[545] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'read'}
    instructions[546] = {5'd1, 4'd2, 4'd4, 16'd5};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'addl'}
    instructions[547] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 15, 'op': 'store'}
    instructions[548] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'literal'}
    instructions[549] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'addl'}
    instructions[550] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'load'}
    instructions[551] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'read'}
    instructions[552] = {5'd1, 4'd2, 4'd4, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'addl'}
    instructions[553] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 16, 'op': 'store'}
    instructions[554] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'literal'}
    instructions[555] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'addl'}
    instructions[556] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'load'}
    instructions[557] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'read'}
    instructions[558] = {5'd0, 4'd2, 4'd0, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'literal': 7, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'literal'}
    instructions[559] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 17, 'op': 'store'}
    instructions[560] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'literal'}
    instructions[561] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'addl'}
    instructions[562] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'load'}
    instructions[563] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'read'}
    instructions[564] = {5'd0, 4'd2, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'literal': 1, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'literal'}
    instructions[565] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 18, 'op': 'store'}
    instructions[566] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'literal'}
    instructions[567] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'addl'}
    instructions[568] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'load'}
    instructions[569] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'read'}
    instructions[570] = {5'd0, 4'd2, 4'd0, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'literal': 6, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'literal'}
    instructions[571] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 19, 'op': 'store'}
    instructions[572] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'literal'}
    instructions[573] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'addl'}
    instructions[574] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'load'}
    instructions[575] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'read'}
    instructions[576] = {5'd1, 4'd2, 4'd4, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'addl'}
    instructions[577] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 20, 'op': 'store'}
    instructions[578] = {5'd0, 4'd8, 4'd0, 16'd14};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'literal': 14, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'literal'}
    instructions[579] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'store'}
    instructions[580] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'addl'}
    instructions[581] = {5'd1, 4'd8, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'addl'}
    instructions[582] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'addl'}
    instructions[583] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'load'}
    instructions[584] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[585] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'load'}
    instructions[586] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'subtract'}
    instructions[587] = {5'd1, 4'd2, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'addl'}
    instructions[588] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 21, 'op': 'store'}
    instructions[589] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'literal'}
    instructions[590] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'store'}
    instructions[591] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'addl'}
    instructions[592] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'literal'}
    instructions[593] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'store'}
    instructions[594] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'addl'}
    instructions[595] = {5'd1, 4'd8, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'addl'}
    instructions[596] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'addl'}
    instructions[597] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'load'}
    instructions[598] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[599] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'load'}
    instructions[600] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'add'}
    instructions[601] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[602] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'load'}
    instructions[603] = {5'd15, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'unsigned_shift_right'}
    instructions[604] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'addl'}
    instructions[605] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 22, 'op': 'store'}
    instructions[606] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'literal'}
    instructions[607] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'store'}
    instructions[608] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[609] = {5'd1, 4'd8, 4'd4, 16'd4};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[610] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[611] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[612] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[613] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[614] = {5'd16, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'equal'}
    instructions[615] = {5'd8, 4'd0, 4'd8, 16'd625};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'label': 625, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[616] = {5'd0, 4'd8, 4'd0, 16'd515};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'literal': 515, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'literal'}
    instructions[617] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'store'}
    instructions[618] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[619] = {5'd1, 4'd8, 4'd4, 16'd5};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[620] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[621] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[622] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[623] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[624] = {5'd16, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'equal'}
    instructions[625] = {5'd8, 4'd0, 4'd8, 16'd635};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'label': 635, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[626] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'literal': 1029, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'literal'}
    instructions[627] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'store'}
    instructions[628] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[629] = {5'd1, 4'd8, 4'd4, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[630] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'addl'}
    instructions[631] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[632] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[633] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'load'}
    instructions[634] = {5'd16, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'equal'}
    instructions[635] = {5'd8, 4'd0, 4'd8, 16'd709};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'a': 8, 'label': 709, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[636] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26, 'op': 'literal'}
    instructions[637] = {5'd1, 4'd2, 4'd4, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26, 'op': 'addl'}
    instructions[638] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 26, 'op': 'store'}
    instructions[639] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27, 'op': 'addl'}
    instructions[640] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27, 'op': 'addl'}
    instructions[641] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27, 'op': 'load'}
    instructions[642] = {5'd8, 4'd0, 4'd8, 16'd698};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 8, 'label': 698, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'jmp_if_false'}
    instructions[643] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'literal'}
    instructions[644] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[645] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[646] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'read'}
    instructions[647] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[648] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[649] = {5'd1, 4'd8, 4'd4, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[650] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[651] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[652] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[653] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[654] = {5'd1, 4'd8, 4'd4, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[655] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[656] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[657] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[658] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[659] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'literal'}
    instructions[660] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[661] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[662] = {5'd1, 4'd8, 4'd4, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[663] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[664] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[665] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[666] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[667] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'add'}
    instructions[668] = {5'd1, 4'd2, 4'd4, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[669] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[670] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[671] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[672] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[673] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[674] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'add'}
    instructions[675] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'addl'}
    instructions[676] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[677] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'load'}
    instructions[678] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 28, 'op': 'store'}
    instructions[679] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[680] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[681] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'load'}
    instructions[682] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'store'}
    instructions[683] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[684] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'literal'}
    instructions[685] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'store'}
    instructions[686] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[687] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[688] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[689] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'load'}
    instructions[690] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[691] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'load'}
    instructions[692] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'subtract'}
    instructions[693] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'addl'}
    instructions[694] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'store'}
    instructions[695] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[696] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 29, 'op': 'load'}
    instructions[697] = {5'd11, 4'd0, 4'd0, 16'd699};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'label': 699, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'goto'}
    instructions[698] = {5'd11, 4'd0, 4'd0, 16'd700};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'label': 700, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'goto'}
    instructions[699] = {5'd11, 4'd0, 4'd0, 16'd639};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27 {'label': 639, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 27, 'op': 'goto'}
    instructions[700] = {5'd1, 4'd8, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'addl'}
    instructions[701] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'addl'}
    instructions[702] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'load'}
    instructions[703] = {5'd0, 4'd2, 4'd0, 16'd4};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'literal': 4, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'literal'}
    instructions[704] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'store'}
    instructions[705] = {5'd1, 4'd3, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'addl'}
    instructions[706] = {5'd1, 4'd4, 4'd7, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'addl'}
    instructions[707] = {5'd12, 4'd0, 4'd6, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31 {'a': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 31, 'op': 'return'}
    instructions[708] = {5'd11, 4'd0, 4'd0, 16'd738};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24 {'label': 738, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 24, 'op': 'goto'}
    instructions[709] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35, 'op': 'addl'}
    instructions[710] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35, 'op': 'addl'}
    instructions[711] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35, 'op': 'load'}
    instructions[712] = {5'd8, 4'd0, 4'd8, 16'd736};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40 {'a': 8, 'label': 736, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40, 'op': 'jmp_if_false'}
    instructions[713] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36, 'op': 'literal'}
    instructions[714] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36, 'op': 'addl'}
    instructions[715] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36, 'op': 'load'}
    instructions[716] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36 {'a': 8, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 36, 'op': 'read'}
    instructions[717] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[718] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[719] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'load'}
    instructions[720] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'store'}
    instructions[721] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[722] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'literal'}
    instructions[723] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'store'}
    instructions[724] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[725] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[726] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[727] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'load'}
    instructions[728] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[729] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'load'}
    instructions[730] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'subtract'}
    instructions[731] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'addl'}
    instructions[732] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'store'}
    instructions[733] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[734] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 37, 'op': 'load'}
    instructions[735] = {5'd11, 4'd0, 4'd0, 16'd737};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40 {'label': 737, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40, 'op': 'goto'}
    instructions[736] = {5'd11, 4'd0, 4'd0, 16'd738};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40 {'label': 738, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 40, 'op': 'goto'}
    instructions[737] = {5'd11, 4'd0, 4'd0, 16'd709};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35 {'label': 709, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 35, 'op': 'goto'}
    instructions[738] = {5'd11, 4'd0, 4'd0, 16'd530};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 12 {'label': 530, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 12, 'op': 'goto'}
    instructions[739] = {5'd1, 4'd3, 4'd3, 16'd3};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45 {'a': 3, 'literal': 3, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45, 'op': 'addl'}
    instructions[740] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'literal'}
    instructions[741] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'store'}
    instructions[742] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'addl'}
    instructions[743] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'literal'}
    instructions[744] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'store'}
    instructions[745] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'addl'}
    instructions[746] = {5'd1, 4'd8, 4'd4, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'addl'}
    instructions[747] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'addl'}
    instructions[748] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'load'}
    instructions[749] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[750] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'load'}
    instructions[751] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'add'}
    instructions[752] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[753] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'load'}
    instructions[754] = {5'd15, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'unsigned_shift_right'}
    instructions[755] = {5'd1, 4'd2, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'addl'}
    instructions[756] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 49, 'op': 'store'}
    instructions[757] = {5'd0, 4'd8, 4'd0, 16'd14};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'literal': 14, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'literal'}
    instructions[758] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'store'}
    instructions[759] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'addl'}
    instructions[760] = {5'd1, 4'd8, 4'd4, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'addl'}
    instructions[761] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'addl'}
    instructions[762] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'load'}
    instructions[763] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[764] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'load'}
    instructions[765] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'add'}
    instructions[766] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'addl'}
    instructions[767] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 50, 'op': 'store'}
    instructions[768] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'literal'}
    instructions[769] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'addl'}
    instructions[770] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'load'}
    instructions[771] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'store'}
    instructions[772] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'addl'}
    instructions[773] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'addl'}
    instructions[774] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'addl'}
    instructions[775] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'load'}
    instructions[776] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[777] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'load'}
    instructions[778] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'write'}
    instructions[779] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 52, 'op': 'addl'}
    instructions[780] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'literal'}
    instructions[781] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'addl'}
    instructions[782] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'load'}
    instructions[783] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'store'}
    instructions[784] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'addl'}
    instructions[785] = {5'd0, 4'd8, 4'd0, 16'd7};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'literal': 7, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'literal'}
    instructions[786] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'addl'}
    instructions[787] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'load'}
    instructions[788] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[789] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'load'}
    instructions[790] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'write'}
    instructions[791] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 53, 'op': 'addl'}
    instructions[792] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'literal'}
    instructions[793] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'addl'}
    instructions[794] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'load'}
    instructions[795] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'store'}
    instructions[796] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'addl'}
    instructions[797] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'literal'}
    instructions[798] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'addl'}
    instructions[799] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'load'}
    instructions[800] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[801] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'load'}
    instructions[802] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'write'}
    instructions[803] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 54, 'op': 'addl'}
    instructions[804] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'literal'}
    instructions[805] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'addl'}
    instructions[806] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'load'}
    instructions[807] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'store'}
    instructions[808] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'addl'}
    instructions[809] = {5'd0, 4'd8, 4'd0, 16'd6};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'literal': 6, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'literal'}
    instructions[810] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'addl'}
    instructions[811] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'load'}
    instructions[812] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[813] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'load'}
    instructions[814] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'write'}
    instructions[815] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 55, 'op': 'addl'}
    instructions[816] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'literal'}
    instructions[817] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'addl'}
    instructions[818] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'load'}
    instructions[819] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'store'}
    instructions[820] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'addl'}
    instructions[821] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'literal'}
    instructions[822] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[823] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'load'}
    instructions[824] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'write'}
    instructions[825] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 56, 'op': 'addl'}
    instructions[826] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'literal'}
    instructions[827] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'addl'}
    instructions[828] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'load'}
    instructions[829] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'store'}
    instructions[830] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'addl'}
    instructions[831] = {5'd0, 4'd8, 4'd0, 16'd515};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'literal': 515, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'literal'}
    instructions[832] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[833] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'load'}
    instructions[834] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'write'}
    instructions[835] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 57, 'op': 'addl'}
    instructions[836] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'literal'}
    instructions[837] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'addl'}
    instructions[838] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'load'}
    instructions[839] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'store'}
    instructions[840] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'addl'}
    instructions[841] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'literal': 1029, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'literal'}
    instructions[842] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[843] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'load'}
    instructions[844] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'write'}
    instructions[845] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 58, 'op': 'addl'}
    instructions[846] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'literal'}
    instructions[847] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'addl'}
    instructions[848] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'load'}
    instructions[849] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'store'}
    instructions[850] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'addl'}
    instructions[851] = {5'd1, 4'd8, 4'd4, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'addl'}
    instructions[852] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'addl'}
    instructions[853] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'load'}
    instructions[854] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[855] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'load'}
    instructions[856] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'write'}
    instructions[857] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 59, 'op': 'addl'}
    instructions[858] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61 {'literal': 0, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61, 'op': 'literal'}
    instructions[859] = {5'd1, 4'd2, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61, 'op': 'addl'}
    instructions[860] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 61, 'op': 'store'}
    instructions[861] = {5'd1, 4'd8, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62, 'op': 'addl'}
    instructions[862] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62, 'op': 'addl'}
    instructions[863] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62, 'op': 'load'}
    instructions[864] = {5'd8, 4'd0, 4'd8, 16'd921};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67 {'a': 8, 'label': 921, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67, 'op': 'jmp_if_false'}
    instructions[865] = {5'd0, 4'd8, 4'd0, 16'd41};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'literal': 41, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'literal'}
    instructions[866] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[867] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[868] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'store'}
    instructions[869] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[870] = {5'd1, 4'd8, 4'd4, -16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[871] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[872] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[873] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'store'}
    instructions[874] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[875] = {5'd1, 4'd8, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[876] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[877] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[878] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'store'}
    instructions[879] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[880] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'literal'}
    instructions[881] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'store'}
    instructions[882] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[883] = {5'd1, 4'd8, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[884] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[885] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[886] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[887] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[888] = {5'd6, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'add'}
    instructions[889] = {5'd1, 4'd2, 4'd4, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[890] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'store'}
    instructions[891] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[892] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[893] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[894] = {5'd5, 4'd2, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[895] = {5'd6, 4'd8, 4'd8, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'add'}
    instructions[896] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[897] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[898] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[899] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'z': 0, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'load'}
    instructions[900] = {5'd13, 4'd0, 4'd0, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 0, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'write'}
    instructions[901] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 63, 'op': 'addl'}
    instructions[902] = {5'd1, 4'd8, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[903] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[904] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'load'}
    instructions[905] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'store'}
    instructions[906] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[907] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'literal': 1, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'literal'}
    instructions[908] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'store'}
    instructions[909] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[910] = {5'd1, 4'd8, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[911] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[912] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 2, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'load'}
    instructions[913] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[914] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'z': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'load'}
    instructions[915] = {5'd10, 4'd8, 4'd8, 16'd10};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'subtract'}
    instructions[916] = {5'd1, 4'd2, 4'd4, 16'd2};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'addl'}
    instructions[917] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 2, 'b': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'store'}
    instructions[918] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'comment': 'pop', 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[919] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64 {'a': 3, 'z': 8, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 64, 'op': 'load'}
    instructions[920] = {5'd11, 4'd0, 4'd0, 16'd922};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67 {'label': 922, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67, 'op': 'goto'}
    instructions[921] = {5'd11, 4'd0, 4'd0, 16'd923};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67 {'label': 923, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 67, 'op': 'goto'}
    instructions[922] = {5'd11, 4'd0, 4'd0, 16'd861};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62 {'label': 861, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 62, 'op': 'goto'}
    instructions[923] = {5'd1, 4'd3, 4'd4, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45, 'op': 'addl'}
    instructions[924] = {5'd1, 4'd4, 4'd7, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45, 'op': 'addl'}
    instructions[925] = {5'd12, 4'd0, 4'd6, 16'd0};///home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45 {'a': 6, 'trace': /home/jon/Projects/Chips-Demo/demo/examples/image_processor/ethernet.h : 45, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //add
        16'd6:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //greater
        16'd7:
        begin
          result <= $signed(operand_a) > $signed(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd8:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //shift_left
        16'd9:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //subtract
        16'd10:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //goto
        16'd11:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //return
        16'd12:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //write
        16'd13:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //read
        16'd14:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //unsigned_shift_right
        16'd15:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //equal
        16'd16:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      2:
      begin
        s_input_eth_in_ack <= 1;
        if (s_input_eth_in_ack && input_eth_in_stb) begin
          result <= input_eth_in;
          write_enable <= 1;
          s_input_eth_in_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_eth_out_stb <= 1;
        s_output_eth_out <= write_value;
        if (output_eth_out_ack && s_output_eth_out_stb) begin
          s_output_eth_out_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_rs232_out_stb <= 1;
        s_output_rs232_out <= write_value;
        if (output_rs232_out_ack && s_output_rs232_out_stb) begin
          s_output_rs232_out_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_in_ack <= 0;
      s_output_eth_out_stb <= 0;
      s_output_rs232_out_stb <= 0;
    end
  end
  assign input_eth_in_ack = s_input_eth_in_ack;
  assign output_eth_out_stb = s_output_eth_out_stb;
  assign output_eth_out = s_output_eth_out;
  assign output_rs232_out_stb = s_output_rs232_out_stb;
  assign output_rs232_out = s_output_rs232_out;

endmodule
